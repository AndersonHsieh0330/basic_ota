** sch_path: /home/andersonhsieh/repo/basic_ota/sky130/pre_layout_sim/nfet_characterization.sch
**.subckt nfet_characterization
XM1 net2 net1 net3 net3 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
V1 net1 net3 0
V2 net2 net3 0.9
**** begin user architecture code


.control
save all @m.xm1.msky130_fd_pr__nfet_01v8[id]
dc V1 0 3 0.01
write nfet_characterization.raw
.endc



** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt

**** end user architecture code
**.ends
.end
